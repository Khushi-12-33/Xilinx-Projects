library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity HADD is
    Port ( A,B : in  STD_LOGIC;
           S,Cout : out  STD_LOGIC);
end HADD;

architecture Behavioral of HADD is

begin


end Behavioral;

